
module	constant	(	 
			  
				   output	logic	[10:0] const1,
					output	logic	[10:0] const2,
					output	logic	[10:0] const3,
					output	logic	[10:0] const4
);

always_comb
begin
	const1 = 32;
	const2 = 32;
	
	const3 = 50;
	const4 = 32;

end
endmodule


